LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY responder IS
PORT(seg7com:OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		seg7data:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		led:OUT STD_LOGIC;
		key1,key2,key3,key4,key5,clk:IN STD_LOGIC
		);
END ENTITY responder;
ARCHITECTURE RTL OF responder IS
COMPONENT EB IS
	PORT(	OP:OUT STD_LOGIC;
			KEY:IN STD_LOGIC;
			CK:IN STD_LOGIC);
END COMPONENT;
SIGNAL ABC:STD_LOGIC_VECTOR(2 DOWNTO 0):="111";
SIGNAL T,ankey5,ankey4,ankey3,ankey2,ankey1,ABCT:STD_LOGIC:='0';
SIGNAL Q,QND,TGB,QC,JFW,BJF:STD_LOGIC:='1';
SHARED VARIABLE QCB,QE,TG:INTEGER RANGE 0 TO 1:=0;
SHARED VARIABLE MODE,WEI,TEAM:INTEGER RANGE 0 TO 4:=0;
SHARED VARIABLE MIN1,MIN2:INTEGER RANGE 0 TO 10:=0;
SHARED VARIABLE numshow,M1,M2,M3,M4:INTEGER RANGE 0 TO 14:=0;
SHARED VARIABLE SEC1,SEC2:INTEGER RANGE 0 TO 69:=0;
SHARED VARIABLE AS,BS,CS:INTEGER RANGE 0 TO 100:=0;
BEGIN
ABC<=ankey1&ankey2&ankey3;
ABCT<=ankey1 AND ankey2 AND ankey3;
led<=NOT Q;
CHANGETIME:PROCESS(ABCT,ABC,TGB,JFW) IS
BEGIN
	IF(ABCT'EVENT AND ABCT='0')THEN
		IF Q='1' THEN
			IF MODE=0 THEN
				CASE ABC IS
					WHEN "110"=>SEC2:=SEC2+1;IF SEC2>59 THEN SEC2:=0;END IF;TG:=1;
					WHEN "101"=>SEC2:=SEC2+10;IF SEC2>59 THEN SEC2:=SEC2 MOD 10;END IF;TG:=1;
					WHEN "011"=>MIN2:=MIN2+1;IF MIN2>9 THEN MIN2:=0;END IF;TG:=1;
					WHEN OTHERS=>NULL;
				END CASE;
			END IF;
		ELSE
			IF QE=0 THEN
				IF QC='1' THEN
					CASE ABC IS
						WHEN "110"=>TEAM:=3;QC<='0';
						WHEN "101"=>TEAM:=2;QC<='0';
						WHEN "011"=>TEAM:=1;QC<='0';
						WHEN OTHERS=>NULL;
					END CASE;
				END IF;
			END IF;
		END IF;
	END IF;
	IF TGB='0'THEN
		TG:=0;
	END IF;
	IF JFW='0'THEN
		QC<='1';
	END IF;
END PROCESS CHANGETIME;
CHANGEMODE:PROCESS(ankey5,JFW) IS
BEGIN
	IF(ankey5'EVENT AND ankey5='1')THEN		
		IF Q='1' THEN
			MODE:=MODE+1;
			IF MODE=4 THEN
				MODE:=0;
			END IF;		
		END IF;
		IF QCB=1 THEN
			BJF<='0';
		END IF;	
	END IF;
	IF JFW='0' THEN
		BJF<='1';
	END IF;
END PROCESS CHANGEMODE;
START:PROCESS(ankey4,QND,QC,BJF)
BEGIN
	IF(ankey4'EVENT AND ankey4='0')THEN
		IF MODE=0 THEN
			IF QCB=1 THEN
				CASE TEAM IS
					WHEN 1=>AS:=AS+1;
					WHEN 2=>BS:=BS+1;
					WHEN 3=>CS:=CS+1;
					WHEN OTHERS=>NULL;
				END CASE;
				JFW<='0';
			ELSE
				Q<='0';
			END IF;
		END IF;
	END IF;
	IF BJF='0' THEN
		JFW<='0';
	END IF;
	IF QC='1' THEN
		JFW<='1';
	END IF;
	IF QND='0' THEN
		Q<='1';
	END IF;
END PROCESS START;
HC7447:PROCESS(T,JFW)
VARIABLE COUNT1 :INTEGER RANGE 0 TO 500;
VARIABLE COUNT2 :INTEGER RANGE 0 TO 500;  
BEGIN
	IF(T'EVENT AND T='1')THEN
		QND<='1';
		TGB<='1';
		COUNT1:=COUNT1+1;
		IF(COUNT1=500)THEN
			IF QE=0 THEN
				IF Q='0' THEN
					IF QC='1' THEN
						IF SEC1=0 THEN
							IF MIN1=0 THEN
								QE:=1;
							ELSE
								MIN1:=MIN1-1;
								SEC1:=59;
							END IF;
						ELSE
							SEC1:=SEC1-1;
						END IF;
					END IF;
				END IF;
			END IF;
			COUNT1:=0;
		END IF;
		IF QE=1 THEN
			M1:=13;M2:=13;M3:=13;M4:=13;
			COUNT2:=COUNT2+1;
			IF(COUNT2=50)THEN		
				QND<='0';
				COUNT2:=0;
				QE:=0;
				SEC1:=SEC2;
				MIN1:=MIN2;
			END IF;
		ELSE
			IF QC='0' THEN
				CASE TEAM IS
					WHEN 1=>M1:=AS REM 10;M2:=AS/10;M3:=13;M4:=10;
					WHEN 2=>M1:=BS REM 10;M2:=BS/10;M3:=13;M4:=11;
					WHEN 3=>M1:=CS REM 10;M2:=CS/10;M3:=13;M4:=12;
					WHEN OTHERS=>NULL;
				END CASE;
				QCB:=1;
			ELSE
				CASE MODE IS
					WHEN 1=>M1:=AS REM 10;M2:=AS/10;M3:=13;M4:=10;
					WHEN 2=>M1:=BS REM 10;M2:=BS/10;M3:=13;M4:=11;
					WHEN 3=>M1:=CS REM 10;M2:=CS/10;M3:=13;M4:=12;
					WHEN 0=>IF TG=1 THEN SEC1:=SEC2;MIN1:=MIN2;TGB<='0';END IF;M1:=SEC1 REM 10;M2:=SEC1/10;M3:=13;M4:=MIN1;		
					WHEN OTHERS=>NULL;
				END CASE;
			END IF;
		END IF;
		CASE WEI IS
			WHEN 0=>seg7com<="0111";numshow:=M1;
			WHEN 1=>seg7com<="1011";numshow:=M2;
			WHEN 2=>seg7com<="1101";numshow:=M3;
			WHEN 3=>seg7com<="1110";numshow:=M4;
			WHEN OTHERS=>seg7com<="1111";
		END CASE;
		WEI:=WEI+1;
		IF WEI=4 THEN
			WEI:=0;
		END IF;
		seg7data<="11111111";
		CASE numshow IS
			WHEN 0=>seg7data<="11000000";
			WHEN 1=>seg7data<="11111001";
			WHEN 2=>seg7data<="10100100";
			WHEN 3=>seg7data<="10110000";
			WHEN 4=>seg7data<="10011001";
			WHEN 5=>seg7data<="10010010";
			WHEN 6=>seg7data<="10000010";
			WHEN 7=>seg7data<="11111000";
			WHEN 8=>seg7data<="10000000";
			WHEN 9=>seg7data<="10010000";
			WHEN 10=>seg7data<="10001000";
			WHEN 11=>seg7data<="10000011";
			WHEN 12=>seg7data<="11000110";
			WHEN 13=>seg7data<="10111111";
			WHEN 14=>seg7data<="11111111";
		END CASE;
	END IF;
	IF JFW='0' THEN
		SEC1:=SEC2;
		MIN1:=MIN2;
		QND<='0';
		QCB:=0;
	END IF;
END PROCESS HC7447;
HZ1k:PROCESS(clk) IS
VARIABLE CNT:INTEGER:=0;
BEGIN
	IF(clk'EVENT AND clk='1')THEN
		CNT:=CNT+1;
		IF CNT=50000 THEN
			T<=NOT T;
			CNT:=0;
		END IF;
	END IF;
END PROCESS HZ1k;
EB1:EB PORT MAP(ankey1,key1,clk);
EB2:EB PORT MAP(ankey2,key2,clk);
EB3:EB PORT MAP(ankey3,key3,clk);
EB4:EB PORT MAP(ankey4,key4,clk);
EB5:EB PORT MAP(ankey5,key5,clk);
END ARCHITECTURE RTL;