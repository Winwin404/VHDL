LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
ENTITY EB IS
PORT(	OP:OUT STD_LOGIC;
		KEY:IN STD_LOGIC;
		CK:IN STD_LOGIC);
END ENTITY EB;
ARCHITECTURE RTL OF EB IS
BEGIN
PROCESS(CK)
	VARIABLE COUT:INTEGER RANGE 0 TO 100000; 
BEGIN 
	IF KEY='0' THEN 
		IF(CK'EVENT AND CK='1')THEN   --shangshengyan
			IF COUT<10000 THEN 
				COUT:=COUT+1; 
			ELSE 
				COUT:=COUT; 
			END IF; 
			IF COUT=9999 THEN 
				OP<='0'; 
			ELSE 
				OP<='1'; 
			END IF; 
		END IF; 
	ELSE 
		COUT:=0;
	END IF; 
END PROCESS;
END ARCHITECTURE RTL;